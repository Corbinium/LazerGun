** Profile: "SCHEMATIC1-laserSight"  [ C:\Users\corbb\Documents\workspace\LazerGun\Circuit\laserGun2-PSpiceFiles\SCHEMATIC1\laserSight.sim ] 

** Creating circuit file "laserSight.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\corbb\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\23.1.0\PSpice.ini file:
.lib "C:\Users\corbb\Documents\School\ECE_2280\HW\customComponents\CD4007.lib" 
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1s 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
